
module control_unit_top(
    input [6:0] opcode,
    input [2:0] funct3,
    input [6:0] funct7,
    output RegWrite,
    output MemToReg,
    output MemRead,
    output MemWrite,
    output [3:0] ALUOp,
    output ALUSrc,
    output RWsel
);

wire [5:0] mapped_address;

// address_mapper
address_mapper addr_mapper (
    .opcode(opcode),
    .funct3(funct3),
    .funct7(funct7),
    .mapped_address(mapped_address)
);

// control_rom
control_rom ctrl_rom (
    .mapped_address(mapped_address),
    .RegWrite(RegWrite),
    .MemToReg(MemToReg),
    .MemRead(MemRead),
    .MemWrite(MemWrite),
    .ALUOp(ALUOp),
    .ALUSrc(ALUSrc),
    .RWsel(RWsel)
);

endmodule
