module ROB(
    input wire clk,                      // Clock signal
    input wire rst,                      // Reset signal
    input wire ROB_Flush,                // ROB Flush signal
    input wire [31:0] IF_ID_instOut,     // Input instruction (expanded to 32 bits)
    input wire reg_write,                // Register write enable signal from the decode stage
    input wire [31:0] PC,                // Current PC value (expanded to 32 bits)
    input wire ID_excpetion,
    
    input wire alu_exec_done,            // ALU execution completion signal
    input wire [31:0] alu_exec_value,    // ALU executed value
    input wire [31:0] alu_exec_PC,       // ALU execution index

    input wire mul_exec_done,            // Multiplier execution completion signal
    input wire [31:0] mul_exec_value,    // Multiplier executed value
    input wire [31:0] mul_exec_PC,       // Multiplier execution index

    input wire div_excpetion,
    input wire div_exec_done,            // Divider execution completion signal
    input wire [31:0] div_exec_value,    // Divider executed value
    input wire [31:0] div_exec_PC,       // Divider execution index
    
    input wire PcSrc,                    // Branch signal (acts like a done signal)
    input wire [31:0] PC_Return,         // Jump address
    input wire [31:0] branch_index,      // Branch index in ROB
    input wire BR_Done,                

    input wire P_Done,
    input wire [31:0] P_Data,
    input wire [31:0] P_inst_num,

    input wire LS_exception,
    input wire Load_Done,
    input wire [31:0] Store_Addr,
    input wire [31:0] Load_Data,
    input wire [31:0] Load_inst_num,
    
    output reg [31:0] out_value,         // Output value
    output reg [4:0] out_dest,           // Output register destination extracted from instr[11:7]
    output reg out_reg_write,            // Output RegWrite signal to indicate a register write operation
    output reg [31:0] out_Addr,
    output reg exception_sig
);

// ROB memory
    reg [99:0] rob_entry [0:63];            // ROB entry: new_bit(1), ready(1), reg_write(1), value(32), instr(32), PC(32)
    reg [31:0] Store_Addrs [0:63];
    reg [5:0] head;                        // Head pointer (5 bits for 32 entries)
    reg [5:0] tail;                        // Tail pointer (5 bits for 32 entries)
    integer i;

// Reset ROB entries
task reset_rob_entries;
    begin
        for (i = 0; i < 64; i = i + 1) begin
            rob_entry[i] <= 100'b0;     // Reset ROB entry with all fields set to 0
            Store_Addrs[i] <= 32'b0;
        end
    end
endtask

// ROB control logic
always @(posedge clk) begin
    if (rst) begin
        head <= 0;
        tail <= 0;
        reset_rob_entries();
    end else begin
        
        if (PcSrc) begin
            // Update the branch entry with PC_Return value
            for (i = 0; i < 64; i = i + 1) begin
                if (rob_entry[i][31:0] == branch_index) begin
                    rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], PC_Return, rob_entry[i][63:32], rob_entry[i][31:0]};
                    tail <= (i + 1) % 64; // Move tail to the entry right after the branch entry
                    rob_entry[(i+1)%64][98:0] <= 0; // Flush under tail entry
                    rob_entry[(i+2)%64][98:0] <= 0; // Fulsh under tail entry
  
                end
            end
        end else if (IF_ID_instOut != 32'b0) begin  // Only increment tail if the instruction is not invalid (i.e., not a bubble)
            if (ID_exception == 1'b0) begin
                rob_entry[tail] <= {1'b0, 1'b1, 1'b0, reg_write, 32'b0, IF_ID_instOut, PC}; // Store input data in the ROB entry with value set to 32'b0 and new_bit set to 1
                tail <= (tail + 1) % 64;                // Circular buffer handling
            end else begin
                exception_sig <= 1'b1;
                head <= 0;
                tail <= 0;
                reset_rob_entries(); 
            end
        end

        
        // Update the value and set ready flag upon execution completion
        
            for (i = 0; i < 64; i = i + 1) begin
                if (rob_entry[i][98]) begin // Check if the new bit is set to 1
                    if ( alu_exec_done &&rob_entry[i][31:0] == alu_exec_PC) begin
                        rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], alu_exec_value, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC
                    end
                    if ( mul_exec_done && rob_entry[i][31:0] == mul_exec_PC) begin
                        rob_entry[i][99:0] <= {rob_entry[i][98], 1'b1, rob_entry[i][96], mul_exec_value, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC       
                    end
                    if ( div_exec_done &&rob_entry[i][31:0] == div_exec_PC) begin
                        if (LS_exception == 1'b1) begin
                            rob_entry[i][99:0] <= {1'b1, rob_entry[i][98], 1'b1, rob_entry[i][96], div_exec_value, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC  
                        end else begin
                            rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], div_exec_value, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC     
                        end
                    end
                    if ( BR_Done&& rob_entry[i][31:0] == branch_index) begin
                        rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], PC_Return, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC
                    end
                    if ( P_Done&& rob_entry[i][31:0] == P_inst_num) begin
                        rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], P_Data, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC
                    end
                    if ( Load_Done&& rob_entry[i][31:0] == Load_inst_num) begin
                        if (LS_exception == 1'b1) begin
                            rob_entry[i][99:0] <= {1'b1, rob_entry[i][98], 1'b1, rob_entry[i][96], Load_Data, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC
                            Store_Addrs[i][31:0] <= Store_Addr;
                        end else begin
                            rob_entry[i][99:0] <= {rob_entry[i][99], rob_entry[i][98], 1'b1, rob_entry[i][96], Load_Data, rob_entry[i][63:32], rob_entry[i][31:0]}; // Update value and maintain new_bit, reg_write, instr, PC
                            Store_Addrs[i][31:0] <= Store_Addr;
                        end
                    end
                end
            end
        
            if (rob_entry[head][97]) begin       // Check if the entry is ready
                if (rob_entry[head][99] == 1'b0) begin
                    out_value <= rob_entry[head][95:64];     // Output value
                    out_dest <= rob_entry[head][43:39];      // Extract out_dest from instr[11:7]
                    out_reg_write <= rob_entry[head][96];   // Output RegWrite status
                    out_Addr <= Store_Addrs[head][31:0];
                    exception_sig <= 1'b0;
                    rob_entry[head] <= 0;            // Clear the ready flag after consuming the entry
                    head <= (head + 1) % 64;                 // Circular buffer handling
                end else begin
                    exception_sig <= 1'b1;
                    head <= 0;
                    tail <= 0;
                    reset_rob_entries();
                end
            end else begin
                    out_value <= 0;     // Output value
                    out_dest <= 0;      // Extract out_dest from instr[11:7]
                    out_reg_write <= 0;   // Output RegWrite status
                    out_Addr <= 32'd1025;
                    exception_sig <= 0;
            end
        
    end
end




endmodule
