module control_rom(
    input [5:0] mapped_address,
    input reset, // �뵳�딅�� 占쎈뻿占쎌깈 �빊遺쏙옙
    output RegWrite,
    output MemToReg,
    output MemRead,
    output MemWrite,
    output [3:0] ALUOp,
    output [1:0] ALUSrc,
    output RWsel,
    output Branch,
    output Jump, // �빊遺쏙옙占쎈쭆 Jump 占쎈뻿占쎌깈
    output mret,
    output ID_exception
);

reg [12:0] ROM [0:63]; // ROM 占쎄쾿疫꿸퀡占쏙옙 13�뜮袁る뱜嚥∽옙 筌앹빓占�

    assign {mret, RegWrite, MemToReg, MemRead, MemWrite, ALUOp, ALUSrc, RWsel, Branch, Jump} = ROM[mapped_address];

    always @(posedge reset) begin
   
        // 筌뤴뫀諭� 占쎌젫占쎈선 占쎈뻿占쎌깈�몴占� 雅뚯눘�꺖 0占쎈퓠占쎄퐣 0占쎌몵嚥∽옙 �룯�뜃由곤옙�넅
        ROM[0] = 14'b0_0_0_0_0_0000_00_0_0_0;

        // R-占쏙옙占쎌뿯 筌뤿굝議딉옙堉�
        ROM[1] = 14'b0_1_0_0_0_0010_10_0_0_0; // ADD
        ROM[2] = 14'b0_1_0_0_0_0110_10_0_0_0; // SUB
        ROM[3] = 14'b0_1_0_0_0_0000_10_0_0_0; // AND
        ROM[4] = 14'b0_1_0_0_0_0001_10_0_0_0; // OR
        ROM[5] = 14'b0_1_0_0_0_0011_10_0_0_0; // XOR
        ROM[6] = 14'b0_1_0_0_0_0100_10_0_0_0; // SLL
        ROM[7] = 14'b0_1_0_0_0_0101_10_0_0_0; // SRL
        ROM[8] = 14'b0_1_0_0_0_0111_10_0_0_0; // SRA
        ROM[9] = 14'b0_1_0_0_0_1000_10_0_0_0; // SLT
        ROM[10] = 14'b0_1_0_0_0_1001_10_0_0_0; // SLTU

        // 嚥≪뮆諭� 獄쏉옙 占쎈뮞占쎈꽅占쎈선
        ROM[11] = 14'b0_1_1_1_0_0010_11_0_0_0; // 嚥≪뮆諭�
        ROM[12] = 14'b0_0_0_0_1_0010_11_0_0_0; // 占쎈뮞占쎈꽅占쎈선

        // Branch 筌뤿굝議딉옙堉�
        ROM[13] = 14'b0_0_0_0_0_0110_10_0_1_0; // �겫袁㏓┛ 筌뤿굝議딉옙堉깍옙肉� 占쏙옙占쎈립 ALUOp 占쎄퐬占쎌젟

        // I-占쏙옙占쎌뿯 筌앸맩�뻻揶쏉옙 占쎈염占쎄텦 獄쏉옙 ALU 筌뤿굝議딉옙堉�
        ROM[14] = 14'b0_1_0_0_0_0010_11_0_0_0; // ADDI
        ROM[15] = 14'b0_1_0_0_0_1000_11_0_0_0; // SLTI
        ROM[16] = 14'b0_1_0_0_0_1001_11_0_0_0; // SLTIU
        ROM[17] = 14'b0_1_0_0_0_0011_11_0_0_0; // XORI
        ROM[18] = 14'b0_1_0_0_0_0001_11_0_0_0; // ORI
        ROM[19] = 14'b0_1_0_0_0_0000_11_0_0_0; // ANDI
        ROM[20] = 14'b0_1_0_0_0_0100_11_0_0_0; // SLLI
        ROM[21] = 14'b0_1_0_0_0_0101_11_0_0_0; // SRLI
        ROM[22] = 14'b0_1_0_0_0_0111_11_0_0_0; // SRAI

        // LUI, AUIPC, JAL, JALR
        ROM[23] = 14'b0_1_0_0_0_0010_11_0_0_0; // LUI
        ROM[24] = 14'b0_1_0_0_0_0010_01_0_0_0; // AUIPC
        ROM[25] = 14'b0_1_0_0_0_0010_01_1_0_1; // JAL
        ROM[26] = 14'b0_1_0_0_0_0010_11_1_0_1; // JALR

        // �빊遺쏙옙占쎈쭆 筌뤿굝議딉옙堉�
        ROM[27] = 14'b0_1_0_0_0_1010_10_0_0_0; // MUL
        ROM[28] = 14'b0_1_0_0_0_0001_10_0_0_0; // DIV (筌륅옙)
        ROM[29] = 14'b0_1_0_0_0_0000_10_0_0_0; // REM (占쎄돌�솒紐꾬옙)
        //csr inst
        ROM[30] = 14'b0_1_0_0_0_0011_10_0_0_0; //csrrw
        ROM[31] = 14'b0_1_0_0_0_0000_10_0_0_0; //csrc
        ROM[32] = 14'b0_1_0_0_0_0001_10_0_0_0; //csrs
        ROM[33] = 14'b0_1_0_0_0_0011_11_0_0_0; //csrrwi
        ROM[34] = 14'b0_1_0_0_0_0001_11_0_0_0; //csrsi
        ROM[35] = 14'b0_1_0_0_0_0000_11_0_0_0; //csrci
        //mret inst
        ROM[36] = 14'b1_0_0_0_0_0011_10_0_0_0; //mret
//0_1_0_0_0_0011_10_0_0_0 csrrw
//0_1_0_0_0_0001_10_0_0_0 csrs
//0_1_0_0_0_0000_10_0_0_0 csrc
//0_1_0_0_0_0011_11_0_0_0 csrrwi
//0_1_0_0_0_0001_11_0_0_0 csrsi
//0_1_0_0_0_0000_11_0_0_0 csrci

//1_0_0_0_0_0011_10_0_0_0 mret
end
    always @(*) begin
        if( mapped_address == 6d'63)
            ID_exception = 1;
        end else begin
            ID_exception = 0;
    end
endmodule
