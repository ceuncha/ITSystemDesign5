module add4(
    input [31:0] in,  // 입력 신호
    output [31:0] out // 출력 신호
);

assign out = in + 4;

endmodule
